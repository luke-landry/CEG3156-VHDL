library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

library altera_mf;
use altera_mf.all;

entity data_mem is
    port (
        address : in std_logic_vector(7 downto 0);
        clock   : in std_logic;
        data    : in std_logic_vector(7 downto 0);
        wren    : in std_logic;
        q       : out std_logic_vector(7 downto 0)
    );
end entity;

architecture rtl of data_mem is
    component altsyncram
        generic (
            operation_mode => string := "SINGLE_PORT",
            width_a        => integer := 8,
            numwords_a     => 256,
            widthad_a      => 8,
            outdata_reg_a  => string := "UNREGISTERED",
            init_file      => string := "data_mem.mif"
        );
        port (
            address_a : in std_logic_vector(7 downto 0);
            clock0    : in std_logic;
            data_a    : in std_logic_vector(7 downto 0);
            wren_a    : in std_logic;
            q_a       : out std_logic_vector(7 downto 0)
        );
    end component;
begin
    ram_inst: altsyncram
        generic map (
            operation_mode => "SINGLE_PORT",
            width_a        => 8,
            numwords_a     => 256,
            widthad_a      => 8,
            outdata_reg_a  => "UNREGISTERED",
            init_file      => "data_mem.mif"
        )
        port map (
            address_a => address,
            clock0    => clock,
            data_a    => data,
            wren_a    => wren,
            q_a       => q
        );
end architecture;
